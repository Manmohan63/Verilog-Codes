module AND_2_dataflow (output Y, input A, B);
	assign Y = A & B; 
endmodule