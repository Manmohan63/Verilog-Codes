module AND_2_gate (output c, input a, b);  
  and (c, a, b);   // c is the output, a and b are inputs 
endmodule 