module hello;
  initial 
    begin
       $display("Hello, World");
	   $write ("Introduction ");
	   $write ("to Verilog ");
	   $display("Hello, World");
	   $write ("Thank You");
      $finish ;
    end
endmodule 