module 4_bit_adder() ();
    
endmodule